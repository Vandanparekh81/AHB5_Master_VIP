class ahb5_slave_dummy_driver;
  logic [31:0] Hrdata;
  logic Hresp;
  logic Hready;
  logic [DATA_WIDTH-1:0] mem [$];
    
