parameter ADDR_WIDTH = 32; // Addr_Width
parameter DATA_WIDTH = 64; // Data_Width
