parameter DATA_WIDTH = 32;
parameter ADDR_WIDTH = 32;
